library verilog;
use verilog.vl_types.all;
entity Adder_Display is
    port(
        \5H6\           : out    vl_logic;
        B0              : in     vl_logic;
        B1              : in     vl_logic;
        B2              : in     vl_logic;
        B3              : in     vl_logic;
        \5H5\           : out    vl_logic;
        \5H3\           : out    vl_logic;
        \5H2\           : out    vl_logic;
        \5H1\           : out    vl_logic;
        \5H0\           : out    vl_logic;
        \5H4\           : out    vl_logic;
        \4H6\           : out    vl_logic;
        \4H5\           : out    vl_logic;
        \4H4\           : out    vl_logic;
        \4H3\           : out    vl_logic;
        \4H2\           : out    vl_logic;
        \4H1\           : out    vl_logic;
        \4H0\           : out    vl_logic;
        \6H0\           : out    vl_logic;
        A0              : in     vl_logic;
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        A3              : in     vl_logic;
        \6H1\           : out    vl_logic;
        \6H2\           : out    vl_logic;
        \6H3\           : out    vl_logic;
        \6H4\           : out    vl_logic;
        \6H5\           : out    vl_logic;
        \6H6\           : out    vl_logic;
        \7H0\           : out    vl_logic;
        \7H1\           : out    vl_logic;
        \7H2\           : out    vl_logic;
        \7H3\           : out    vl_logic;
        \7H4\           : out    vl_logic;
        \7H5\           : out    vl_logic;
        \7H6\           : out    vl_logic;
        \0H0\           : out    vl_logic;
        \0H1\           : out    vl_logic;
        \0H2\           : out    vl_logic;
        \0H3\           : out    vl_logic;
        \0H4\           : out    vl_logic;
        \0H5\           : out    vl_logic;
        \0H6\           : out    vl_logic;
        \1H0\           : out    vl_logic;
        \1H1\           : out    vl_logic;
        \1H2\           : out    vl_logic;
        \1H3\           : out    vl_logic;
        \1H4\           : out    vl_logic;
        \1H5\           : out    vl_logic;
        \1H6\           : out    vl_logic;
        Q0              : out    vl_logic;
        Q1              : out    vl_logic;
        Q2              : out    vl_logic;
        Q3              : out    vl_logic;
        LED             : out    vl_logic
    );
end Adder_Display;
